

module vga_top(input logic        clk,
	        input logic 	   reset,
		input logic [15:0]  writedata,
		input logic 	   write,
		input 		   chipselect,
		input logic [2:0]  address,
    
    output logic [15:0] readdata,
		output logic [7:0] VGA_R, VGA_G, VGA_B,
		output logic 	   VGA_CLK, VGA_HS, VGA_VS,
		                   VGA_BLANK_n,
		output logic 	   VGA_SYNC_n);

// current VGA pixel coord
   logic [10:0]	   hcount;
   logic [9:0]     vcount;

   logic [7:0] 	   background_r, background_g, background_b;
   logic [15:0]  hv_count;

   parameter BALL_SIZE = 64; // ball size = 64 * 64 pixels

  // actual effective coord to draw ball.
   logic [10:0] ball_x_eff;
   logic [9:0] ball_y_eff;
	
  // pending to update ball's coord (from sw)
  logic [10:0] ball_x_pend;
  logic [9:0] ball_y_pend;

  logic ball_update_pending, ball_x_update_pending, ball_y_update_pending;
  
  assign ball_update_pending = ball_x_update_pending & ball_y_update_pending;

   vga_counters counters(.clk50(clk), .*);

   always_ff @(posedge clk) begin
     if (reset) begin
	background_r <= 8'h0;
	background_g <= 8'h0;
	background_b <= 8'h80;
  ball_x_eff <= 11'd100;  // default
  ball_y_eff <= 10'd100;  // default
  ball_x_pend <= 11'd100;
  ball_y_pend <= 10'd100;
  ball_x_update_pending<= 1'b0;
  ball_y_update_pending<= 1'b0;
  end else begin 
    if (chipselect) begin
      if (write) begin
       case (address)
	 3'h0 : background_r <= writedata[7:0];
	 3'h1 : background_g <= writedata[7:0];
	 3'h2 : background_b <= writedata[7:0];
   3'h3: begin
          ball_x_pend <= writedata[10:0];
          ball_x_update_pending<= 1'b1;
        end
  3'h4: begin
          ball_y_pend <= writedata[9:0];
          ball_y_update_pending<= 1'b1;
        end
       endcase
      end  else begin // read
        case (address)
  3'h5 : hv_count <= {5'b0, hcount};
  3'h6 : hv_count <= {6'b0, vcount};
        endcase 
      end
    end

    if ( (vcount[9] | (vcount[8:5] == 4'b1111)) && ball_update_pending) begin
      ball_x_eff <= ball_x_pend;
      ball_x_update_pending <= 1'b0;
      
      ball_y_eff <= ball_y_pend;
      ball_y_update_pending <= 1'b0;
      end
    end
  end

  assign readdata = hv_count;

   always_comb begin
       {VGA_R, VGA_G, VGA_B} = 24'h000000;
       if (VGA_BLANK_n) begin
          logic signed [11:0] dx, dy;
           dx = (hcount >> 1) - (ball_x_eff[10:1] + BALL_SIZE/2);
           dy = vcount - (ball_y_eff + BALL_SIZE/2);
    
           if ((dx*dx + dy*dy) <= ((BALL_SIZE/2)*(BALL_SIZE/2)))
               {VGA_R, VGA_G, VGA_B} = 24'hffffff;
           else
               {VGA_R, VGA_G, VGA_B} = {background_r, background_g, background_b};
       end
   end
	       
endmodule

module vga_counters(
 input logic 	     clk50, reset,
 output logic [10:0] hcount,  // hcount[10:1] is pixel column
 output logic [9:0]  vcount,  // vcount[9:0] is pixel row
 output logic 	     VGA_CLK, VGA_HS, VGA_VS, VGA_BLANK_n, VGA_SYNC_n);

/*
 * 640 X 480 VGA timing for a 50 MHz clock: one pixel every other cycle
 * 
 * HCOUNT 1599 0             1279       1599 0
 *             _______________              ________
 * ___________|    Video      |____________|  Video
 * 
 * 
 * |SYNC| BP |<-- HACTIVE -->|FP|SYNC| BP |<-- HACTIVE
 *       _______________________      _____________
 * |____|       VGA_HS          |____|
 */
   // Parameters for hcount
   parameter HACTIVE      = 11'd 1280,
             HFRONT_PORCH = 11'd 32,
             HSYNC        = 11'd 192,
             HBACK_PORCH  = 11'd 96,   
             HTOTAL       = HACTIVE + HFRONT_PORCH + HSYNC +
                            HBACK_PORCH; // 1600
   
   // Parameters for vcount
   parameter VACTIVE      = 10'd 480,
             VFRONT_PORCH = 10'd 10,
             VSYNC        = 10'd 2,
             VBACK_PORCH  = 10'd 33,
             VTOTAL       = VACTIVE + VFRONT_PORCH + VSYNC +
                            VBACK_PORCH; // 525

   logic endOfLine;
   
   always_ff @(posedge clk50 or posedge reset)
     if (reset)          hcount <= 0;
     else if (endOfLine) hcount <= 0;
     else  	         hcount <= hcount + 11'd 1;

   assign endOfLine = hcount == HTOTAL - 1;
       
   logic endOfField;
   
   always_ff @(posedge clk50 or posedge reset)
     if (reset)          vcount <= 0;
     else if (endOfLine)
       if (endOfField)   vcount <= 0;
       else              vcount <= vcount + 10'd 1;

   assign endOfField = vcount == VTOTAL - 1;

   // Horizontal sync: from 0x520 to 0x5DF (0x57F)
   // 101 0010 0000 to 101 1101 1111
   assign VGA_HS = !( (hcount[10:8] == 3'b101) &
		      !(hcount[7:5] == 3'b111));
   assign VGA_VS = !( vcount[9:1] == (VACTIVE + VFRONT_PORCH) / 2);

   assign VGA_SYNC_n = 1'b0; // For putting sync on the green signal; unused
   
   // Horizontal active: 0 to 1279     Vertical active: 0 to 479
   // 101 0000 0000  1280	       01 1110 0000  480
   // 110 0011 1111  1599	       10 0000 1100  524
   assign VGA_BLANK_n = !( hcount[10] & (hcount[9] | hcount[8]) ) &
			!( vcount[9] | (vcount[8:5] == 4'b1111) );

   /* VGA_CLK is 25 MHz
    *             __    __    __
    * clk50    __|  |__|  |__|
    *        
    *             _____       __
    * hcount[0]__|     |_____|
    */
   assign VGA_CLK = hcount[0]; // 25 MHz clock: rising edge sensitive
   
endmodule
